//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux_2_1
(
  input  [3:0] d0, d1,
  input        sel, // select - выбирает, какой сигнал подать на выход
					// Поскольку 2 входных сигнала, sel однобитный
  output [3:0] y    // По умолчанию тип wire
);

  // тернарный оператор
  // если sel = 1 выбирает d1, иначе d0
  assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module mux_4_1
(
  input  [3:0] d0, d1, d2, d3,
  input  [1:0] sel, // sel двухбитный 11, так как 4 сигнала. 
  output [3:0] y
);

  // Task:
  // Using code for mux_2_1 as an example,
  // write code for 4:1 mux using "?:" operator

	// если первый бит 1, то выбирает между 3 (11) и 2 (10) в зависимости от того, какой второй бит
	// иначе выбирает между 1 (01) и 0 (00)
	assign y = sel[1] ? (sel[0] ? d3 : d2) : (sel[0] ? d1 : d0);


endmodule
