//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux_2_1
(
  input        [3:0] d0, d1,
  input              sel,
  output logic [3:0] y
);

  always_comb
    case (sel)
      1'd0: y = d0;
      1'd1: y = d1;
    endcase

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module mux_4_1
(
  input        [3:0] d0, d1, d2, d3,
  input        [1:0] sel,
  output logic [3:0] y
);

  // Task:
  // Using code for mux_2_1 as an example,
  // write code for 4:1 mux using the "case" statement
  
    // То же самое, что и в предыдущем задании
    // Нужно перебрать все варианты, только теперь через case

    // always_comb блок будет пересчитываться каждый раз, когда изменятеся
    // хотя был один из сигналов внутри него. То есть на y будет всегда подаваться актуальная информация
    always_comb
        case (sel)
        2'b00: y = d0; // Если sel = 00, выход y = d0
        2'b01: y = d1; // Если sel = 01, выход y = d1
        2'b10: y = d2; // Если sel = 10, выход y = d2
        2'b11: y = d3; // Если sel = 11, выход y = d3
        endcase


endmodule
