//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux_4_1_width_2
(
  // Мультиплексор обрабатывает только 2 битные сигналы
  input  [1:0] d0, d1, d2, d3,
  input  [1:0] sel,
  output [1:0] y
);


// Это решение 1 задания
// только тут оно немного другое 
  assign y = sel [1] ? (sel [0] ? d3 : d2)
                     : (sel [0] ? d1 : d0);

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module mux_4_1
(
  // 4 битные сигналы
  input  [3:0] d0, d1, d2, d3,
  input  [1:0] sel,
  output [3:0] y
);

  // Task:
  // Implement mux_4_1 with 4-bit data
  // using two instances of mux_4_1_width_2 with 2-bit data
   

   // Суть задания в том, что у нас есть 4 битные сигналы
   // Но наш мультиплексор обрабатывает только 2 бита

    // Решение состоит в том, что мы разобьём 4 битный сигнал на
    // два 2 битных, каждый из которых обработаем мультиплексором.
    // Затем два 2 битных сигнала соединим в один 4 битный

    // Хранение частей 4 битного сигнала
    wire [1:0] y_10;  
    wire [1:0] y_32; 


    // Обработка двух частоей сигнала
    mux_4_1_width_2 mux_10 (
        .d0(d0[1:0]), 
        .d1(d1[1:0]), 
        .d2(d2[1:0]), 
        .d3(d3[1:0]), 
        .sel(sel),    
        .y(y_10)     
        );

    mux_4_1_width_2 mux_32 (
        .d0(d0[3:2]), 
        .d1(d1[3:2]), 
        .d2(d2[3:2]), 
        .d3(d3[3:2]), 
        .sel(sel),    
        .y(y_32)    
        );

    // конкатенация в один сигнал
    assign y = {y_32, y_10}; // { [3:2], [1:0] }



endmodule
