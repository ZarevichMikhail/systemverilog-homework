//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux_2_1
(
  input  [3:0] d0, d1,
  input        sel,
  output [3:0] y
);

  assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module mux_4_1
(
  input  [3:0] d0, d1, d2, d3,
  input  [1:0] sel,
  output [3:0] y
);

  // Task:
  // Implement mux_4_1 using three instances of mux_2_1

    // Мультиплексор 4 в 1 создадим на основе трёх мультиплексоров 2 в 1.
    // Подадим на два 2 в 1 мультиплексора четыре сигнала. 
    // Получим два выхоодных сигнала,
    // которые передадим в третий мультиплексор


    // Выходы первого и второго мультиплексора. 
    wire [3:0] y_01;
    wire [3:0] y_23;


    // Тут идёт создание экземпляра модуля, созданного ранее
    // 
    // sel[0] Выбирает между 0 и 1, и между 2 и 3
    // и присваеват значения в y_01 и y_23
    mux_2_1 mux_01 (.d0(d0), .d1(d1), .sel(sel[0]), .y(y_01));
    mux_2_1 mux_23 (.d0(d2), .d1(d3), .sel(sel[0]), .y(y_23));


    // Третий мультиплексор
    // На него подаются результаты первых двух
    // sel[1] выбирает между предыдущими результатами 
    mux_2_1 completed_mux(.d0(y_01), .d1(y_23), .sel(sel[1]), .y(y));




endmodule
