//----------------------------------------------------------------------------
// Example
//----------------------------------------------------------------------------

module mux
(
  input  d0, d1,
  input  sel,
  output y
);

  assign y = sel ? d1 : d0;

endmodule

//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module and_gate_using_mux
(
    input  a,
    input  b,
    output o
);

  // Task:
  // Implement and gate using instance(s) of mux,
  // constants 0 and 1, and wire connections

    // Таблица истинности для "И"
    // a b a&b
    // 0 0 0
    // 0 1 0
    // 1 0 0
    // 1 1 1

    // Это можно интерпретировать так:
    // a будет управляющим сигналом
    // Если а = 0, то на выходе всегда 0
    // Если a = 1, то на выходе b

    mux and_gate (
        .d0(1'b0),  // если a = 0, то выводим 0
        .d1(b),     // если a = 1, то выводим b
        .sel(a),    // на sel подаём a
        .y(o)       // 
    );



endmodule
